//
// Global Definitions for the DiRT library.
//
`timescale 1ns/1ps

// Booleans
`define FALSE 1'b0
`define TRUE 1'b1

