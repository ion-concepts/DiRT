//-----------------------------------------------------------------------------
// File:    drat2eth_framer.sv
//
// Author:  Ian Buckley, Ion Concepts LLC.
//
// Description:
// Takes raw DRaT packets as input.
// Encapsulates them as Ethernet/IPv4/UDP.
// Ethernet MAC fields and IPv4 address fields are set from CSR's and global for all packet flows.
//
// This module supports 2 methods to map FlowID.DST to UDP Ports.
// If FlowID.DST[8] is set then csr_udp_dst8 sets the upper 10bits of UDP DST port
// and flowID.DST[5:0] set the lower 6 bits.
// If FlowID.DST[8] is clear then flowID.DST[2:0] select from csr_udp_dst[0:7]
// to fully map FlowID.DST top an arbitrary UDP port.
//
// Many header fields are hard coded as local params to sensible value,
// and UDP checksum generation is dissabled.
//
// License: CERN-OHL-P (See LICENSE.md)
//
//-----------------------------------------------------------------------------
`include "global_defs.svh"
`include "ethernet.sv"
`include "drat_protocol.sv"
module drat2eth_framer
  (

   input logic        clk,
   input logic        rst,
   // CSR interface
   input logic [47:0] csr_mac_dst,
   input logic [47:0] csr_mac_src,
   input logic [31:0] csr_ipv4_dst,
   input logic [31:0] csr_ipv4_src,
   input logic [15:0] csr_udp_src,
   input logic [15:0] csr_udp_dst0,
   input logic [15:0] csr_udp_dst1,
   input logic [15:0] csr_udp_dst2,
   input logic [15:0] csr_udp_dst3,
   input logic [15:0] csr_udp_dst4,
   input logic [15:0] csr_udp_dst5,
   input logic [15:0] csr_udp_dst6,
   input logic [15:0] csr_udp_dst7,
   input logic [9:0]  csr_udp_dst8,


   input logic        csr_enable,
   output logic       csr_idle,
   // DRaT protocol input bus (64b TDATA)
   axis_t.slave in_axis,
   // Ethernet/IPv4/UDP encapsulated output bus (68b TDATA)
   axis_t.master out_axis

   );

   // Constants
   localparam logic [15:0] C_ETHERTYPE = 16'h0800;
   localparam logic [3:0]  C_VERSION = 4'd4;         // IPv4
   localparam logic [3:0]  C_IHL = 4'd5;             // Standard IPv4 header with no options
   localparam logic [7:0]  C_DSCP_ECN = 8'd0;        // DSCP and ECN unused
   localparam logic [15:0] C_IDENTIFICATION = 16'd0; // Unused
   localparam logic [2:0]  C_FLAGS = 3'b010;         // Don't fragment
   localparam logic [12:0] C_FRAGMENT_OFFSET = 13'd0;// Don't fragment
   localparam logic [7:0]  C_TIME_TO_LIVE = 8'd16;   // TTL
   localparam logic [7:0]  C_PROTOCOL = 8'd17;       // UDP
   localparam logic [15:0] C_UDP_CHECKSUM = 16'd0;   // UDP checksum dissabled.
   // Precalculate constant parts of IPv4 header checksum
   localparam logic [17:0] C_PRECALC_CHECKSUM = {C_VERSION, C_IHL, C_DSCP_ECN} + {C_FLAGS, C_FRAGMENT_OFFSET} + {C_TIME_TO_LIVE, C_PROTOCOL};


   drat_protocol::pkt_header_t drat_header;
   logic [15:0]            calc_length;
   logic [15:0]            udp_src, udp_dst;
   logic [18:0]            checksum_ipaddr;
   logic [18:0]            checksum_ipaddr_plus_len;
   logic [16:0]            checksum_pre;
   logic [15:0]            ipv4_checksum;


   //-----------------------------------------------------------------------------
   // State machine
   //-----------------------------------------------------------------------------
   enum {
         S_IDLE,
         S_HEADER1,
         S_HEADER2,
         S_HEADER3,
         S_HEADER4,
         S_HEADER5,
         S_HEADER6,
         S_PAYLOAD,
         S_LAST
         } state;

   always_ff @(posedge clk) begin
        if (rst) begin
           state <= S_IDLE;
           drat_header <= '0;
           csr_idle <= 1'b0;

        end else begin
           case (state)
             // Use first beat of new packet to populate DRaT header structure
             S_IDLE: begin
                // Wait for the next DRaT packet to be valid
                if (csr_enable && in_axis.tvalid) begin
                   // Grab DRaT header
                   drat_header <= drat_protocol::populate_header_no_timestamp(in_axis.tdata);
                   state <= S_HEADER1;
                end
                csr_idle <= ~csr_enable;
             end
             // 1st beat of header (Ethernet)
             S_HEADER1: begin
                if (out_axis.tready == 1)
	          state <= S_HEADER2;
             end
             // 2nd beat of header( Ethernet)
             S_HEADER2: begin
               if (out_axis.tready == 1)
	          state <= S_HEADER3;
             end
             // 3rd beat of header (Ethernet/IPv4)
             S_HEADER3: begin
               if (out_axis.tready == 1)
	          state <= S_HEADER4;
             end
             // 4th beat of header (IPv4)
             S_HEADER4: begin
               if (out_axis.tready == 1)
	          state <= S_HEADER5;
             end
             // 5th beat of header (IPv4)
             S_HEADER5: begin
                if (out_axis.tready == 1)
	          state <= S_HEADER6;
            end
             // 6th beat of header (UDP)
             S_HEADER6: begin
               if (out_axis.tready == 1)
	          state <= S_PAYLOAD;
             end
             // subsequent beats of packet
             S_PAYLOAD: begin
                if ((in_axis.tvalid == 1) && (out_axis.tready == 1) && (in_axis.tlast == 1))
	            state <= S_IDLE;
             end
             // Should never get to default
             default: begin
                state <= S_IDLE;
             end
           endcase // case (state)

        end // else: !if(rst)
   end // always_ff @ (posedge clk)

   // Recaclulate IPv4 and UDP packet lengths on the fly to re-use one adder and register.
   always_ff @(posedge clk) begin
      if (rst) begin
         calc_length <= 16'h0;
      end else if (state == S_HEADER1) begin
         calc_length <= drat_header.length + 16'd28;
      end else if (state == S_HEADER4) begin
         calc_length <= drat_header.length + 16'd8;
      end
   end

   // Use 3 LSB's of DRaT Flow_ID to choose from 8 UDP src+dst port tuples (Where src is constant)
   always_comb begin
      // UDP Source is always the same.
      udp_src = csr_udp_src;
      // if FlowID.dst[8] is set we use direct DRat->UDP port map mode.
      if (drat_header.flow_id[8] == 1) begin
         // Direct Map FlowID.dst[5:0] to UDP Port LSBs.
         // csr_udp_dst8 sets 10MSB's of UDP port
         udp_dst = {csr_udp_dst8,drat_header.flow_id[5:0]};
      end else begin
         // Map FlowID.dst[2:0] to individual UDP ports from CSR's
         case(drat_header.flow_id[2:0])
           0: begin
              udp_dst = csr_udp_dst0;
           end
           1:begin
              udp_dst = csr_udp_dst1;
           end
           2:begin
              udp_dst = csr_udp_dst2;
           end
           3:begin
              udp_dst = csr_udp_dst3;
           end
           4: begin
              udp_dst = csr_udp_dst4;
           end
           5:begin
              udp_dst = csr_udp_dst5;
           end
           6:begin
              udp_dst = csr_udp_dst6;
           end
           7:begin
              udp_dst = csr_udp_dst7;
           end
         endcase // case (drat_header.flow_id[2:0])
      end
   end // always_comb


   // AXIS handshaking. These are all Async timing paths through the block
   always_comb begin
      in_axis.tready = (state == S_PAYLOAD) ? out_axis.tready : 1'b0;
      out_axis.tvalid = (state == S_PAYLOAD) ? in_axis.tvalid :  (state == S_IDLE) ? 1'b0 : 1'b1;
      out_axis.tlast = (state == S_PAYLOAD) ? in_axis.tlast : 1'b0;
      out_axis.tdata[67:64] = ((state == S_PAYLOAD) & in_axis.tlast) ? {1'b0,drat_header.length[2:0]} : 4'b0000;
   end

   // Abreviated IPv4 header checksum calc because many fields are constant or pre-programmed.
   // Gate updates with state to capture correct IPv4 length value, fold in carrys out the MSBs, and pipeline for clock speed.
   always_ff @(posedge clk) begin
      if (state == S_HEADER1)
        checksum_ipaddr[18:0] <= csr_ipv4_src[15:0] +  csr_ipv4_dst[15:0] + csr_ipv4_src[31:16] +  csr_ipv4_dst[31:16] + C_PRECALC_CHECKSUM;
      // Add in packet length then fold in 3 bits of carry
      if (state == S_HEADER2)
        checksum_pre[16:0] <= (checksum_ipaddr_plus_len[15:0] + checksum_ipaddr_plus_len[18:16]);
      // Possibility of one more carry bit that needs to fold in
      if (state == S_HEADER3)
        ipv4_checksum[15:0] <= ~(checksum_pre[15:0] + checksum_pre[16]);
   end

   // Enough remaining dynamic range in checksum_ipaddr to add in another 16 bits without generating a carry into [19]
   always_comb begin
      checksum_ipaddr_plus_len[18:0] = checksum_ipaddr[18:0] + calc_length[15:0];
   end

   // Mux TDATA source for egress to inject header fields before payload beats.
   always_comb begin
      case(state)
        S_HEADER1 : out_axis.tdata[63:0] <= { 48'h0, csr_mac_dst[47:32]};
        S_HEADER2 : out_axis.tdata[63:0] <= { csr_mac_dst[31:0], csr_mac_src[47:16]};
        S_HEADER3 : out_axis.tdata[63:0] <= { csr_mac_src[15:0], C_ETHERTYPE, C_VERSION, C_IHL, C_DSCP_ECN, calc_length };
        S_HEADER4 : out_axis.tdata[63:0] <= { C_IDENTIFICATION , C_FLAGS, C_FRAGMENT_OFFSET, C_TIME_TO_LIVE, C_PROTOCOL, ipv4_checksum};
        S_HEADER5 : out_axis.tdata[63:0] <= { csr_ipv4_src, csr_ipv4_dst};
        S_HEADER6 : out_axis.tdata[63:0] <= { udp_src, udp_dst, calc_length, C_UDP_CHECKSUM};
        default : out_axis.tdata[63:0] <= in_axis.tdata[63:0]; // Pass through payload.
      endcase // case (state)
   end

endmodule // drat2eth_framer
