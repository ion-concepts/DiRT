//-------------------------------------------------------------------------------
// File:   global_defs.svh
//
// Author:  Ian Buckley, Ion Concepts LLC
//
// Global Definitions for the DiRT library.
//
//  License: CERN-OHL-P (See LICENSE.md)
//
//-------------------------------------------------------------------------------
`timescale 1ns/1ps

// Booleans
`define FALSE 1'b0
`define TRUE 1'b1

